library verilog;
use verilog.vl_types.all;
entity tbff is
end tbff;
