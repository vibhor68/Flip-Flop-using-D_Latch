library verilog;
use verilog.vl_types.all;
entity tbff2 is
end tbff2;
